//-----------------------------------------------------------------------------
// Title         : Display LUT
// Project       : Clock
//-----------------------------------------------------------------------------
// File          : disp_lut.sv
// Author        : Daniel Sun  <dcsun88osh@gmail.com>
// Created       : 31.10.2018
// Last modified : 31.10.2018
//-----------------------------------------------------------------------------
// Description : Display controller look up table
// 
//-----------------------------------------------------------------------------
// Copyright (c) 2018 by  This model is the confidential and
// proprietary property of  and the possession or use of this
// file requires a written license from .
//------------------------------------------------------------------------------
// Modification history :
// 31.10.2018 : created
//-----------------------------------------------------------------------------

// `begin_keywords "1800-2012"
// `timescale 1ps/1ps

module disp_lut
//  import util_pkg::*;
   (
    input logic         rst_n,
    input logic         clk,

    input logic [9:0]   sram_addr,
    input logic         sram_we,
    input logic [31:0]  sram_datao,
    output logic [31:0] sram_datai,

    input logic [11:0]  lut_addr,
    output logic [7:0]  lut_data
    );


   logic                rst;

   assign rst = ~rst_n;


   // BRAM_TDP_MACRO: True Dual Port RAM
   //                 Virtex-7
   // Xilinx HDL Language Template, version 2014.4
   
   //////////////////////////////////////////////////////////////////////////
   // DATA_WIDTH_A/B | BRAM_SIZE | RAM Depth | ADDRA/B Width | WEA/B Width //
   // ===============|===========|===========|===============|=============//
   //     19-36      |  "36Kb"   |    1024   |    10-bit     |    4-bit    //
   //     10-18      |  "36Kb"   |    2048   |    11-bit     |    2-bit    //
   //     10-18      |  "18Kb"   |    1024   |    10-bit     |    2-bit    //
   //      5-9       |  "36Kb"   |    4096   |    12-bit     |    1-bit    //
   //      5-9       |  "18Kb"   |    2048   |    11-bit     |    1-bit    //
   //      3-4       |  "36Kb"   |    8192   |    13-bit     |    1-bit    //
   //      3-4       |  "18Kb"   |    4096   |    12-bit     |    1-bit    //
   //        2       |  "36Kb"   |   16384   |    14-bit     |    1-bit    //
   //        2       |  "18Kb"   |    8192   |    13-bit     |    1-bit    //
   //        1       |  "36Kb"   |   32768   |    15-bit     |    1-bit    //
   //        1       |  "18Kb"   |   16384   |    14-bit     |    1-bit    //
   //////////////////////////////////////////////////////////////////////////

   BRAM_TDP_MACRO #(
      .BRAM_SIZE("36Kb"), // Target BRAM: "18Kb" or "36Kb" 
      .DEVICE("7SERIES"), // Target device: "7SERIES" 
      .DOA_REG(0),        // Optional port A output register (0 or 1)
      .DOB_REG(0),        // Optional port B output register (0 or 1)
      .INIT_A(36'h00000000), // Initial values on port A output port
      .INIT_B(36'h00000000), // Initial values on port B output port
      .INIT_FILE ("NONE"),
      .READ_WIDTH_A (32),  // Valid values are 1-36 (19-36 only valid when BRAM_SIZE="36Kb")
      .READ_WIDTH_B (8),   // Valid values are 1-36 (19-36 only valid when BRAM_SIZE="36Kb")
      .SIM_COLLISION_CHECK ("ALL"), // Collision check enable "ALL", "WARNING_ONLY", 
                                    //   "GENERATE_X_ONLY" or "NONE" 
      .SRVAL_A(36'h00000000), // Set/Reset value for port A output
      .SRVAL_B(36'h00000000), // Set/Reset value for port B output
      .WRITE_MODE_A("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE" 
      .WRITE_MODE_B("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE" 
      .WRITE_WIDTH_A(32), // Valid values are 1-36 (19-36 only valid when BRAM_SIZE="36Kb")
      .WRITE_WIDTH_B(8),  // Valid values are 1-36 (19-36 only valid when BRAM_SIZE="36Kb")
      .INIT_00(256'h000000000000000000000064006300530075006e00380038002000470050004c),
      .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_02(256'h00220023002400250026002700280029002a002b002c002d002e002f00300031),
      .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000200021),
      .INIT_04(256'h003400350036003700380039003a003b003c003d003e003f0040004100420043),
      .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000320033),
      .INIT_06(256'h0046004700480049004a004b004c004d004e004f005000510052005300540055),
      .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000440045),
      .INIT_08(256'h00580059005a005b005c005d005e005f00600061006200630064006500660067),
      .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000560057),
      .INIT_0A(256'h006a006b006c006d006e006f0070007100720073007400750076007700780079),
      .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000680069),
      .INIT_0C(256'h007c007d007e007f002000200020002000200020002000200020002000200020),
      .INIT_0D(256'h00000000000000000000000000000000000000000000000000000000007a007b),
      .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_10(256'h0020002000200020002000880087002000860085002000840183008200810080),
      .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000200020),
      .INIT_12(256'h0020002000200020008800870020008600850020008401830082008100800020),
      .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000200020),
      .INIT_14(256'h0020002000200088008700200086008500200084018300820081008000200020),
      .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000200020),
      .INIT_16(256'h0020002000880087002000860085002000840183008200810080002000200020),
      .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000200020),
      .INIT_18(256'h0020008800870020008600850020008401830082008100800020002000200020),
      .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000200020),
      .INIT_1A(256'h0088008700200086008500200084018300820081008000200020002000200020),
      .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000200020),
      .INIT_1C(256'h0087002000860085002000840183008200810080002000200020002000200020),
      .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000200088),
      .INIT_1E(256'h0020008600850020008401830082008100800020002000200020002000200020),
      .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000880087),
      .INIT_20(256'h0086008500200084018300820081008000200020002000200020002000200088),
      .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000870020),
      .INIT_22(256'h0085002000840183008200810080002000200020002000200020002000880087),
      .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000200086),
      .INIT_24(256'h0020008401830082008100800020002000200020002000200020008800870020),
      .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000860085),
      .INIT_26(256'h0084018300820081008000200020002000200020002000200088008700200086),
      .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000850020),
      .INIT_28(256'h0183008200810080002000200020002000200020002000880087002000860085),
      .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000200084),
      .INIT_2A(256'h0082008100800020002000200020002000200020008800870020008600850020),
      .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000840183),
      .INIT_2C(256'h0081008000200020002000200020002000200088008700200086008500200084),
      .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000001830082),
      .INIT_2E(256'h0080002000200020002000200020002000880087002000860085002000840183),
      .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000820081),
      .INIT_30(256'h0020002000200020002000200020008800870020008600850020008401830082),
      .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000810080),
      .INIT_32(256'h0020002000200020002000200088008700200086008500200084018300820081),
      .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000800020),
      .INIT_34(256'h002000470050004c002000470050004c002000470050004c002000470050004c),
      .INIT_35(256'h002000470050004c002000470050004c002000470050004c002000470050004c),
      .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_38(256'h000000000000000000000064006300530075006e00380038002000470050004c),
      .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3C(256'h0020008800870020008600850020008401830082008100800020002000200020),
      .INIT_3D(256'h0020002000200020002000200020002000200020002000200020002000200020),
      .INIT_3E(256'h0138013801380138013801380138013801380138013801380138013801380138),
      .INIT_3F(256'h0138013801380138013801380138013801380138013801380138013801380138),
      
      // The next set of INIT_xx are valid when configured as 36Kb
      .INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_41(256'hca0012000000f6fee0beb666f2da60fc00010200000000000400000000440000),
      .INIT_42(256'h1000000000da766e547c7c1eb6ccd6cefceca81cae780c6ebc8e9e7a9cfeee00),
      .INIT_43(256'h0080000000da766e4438381eb60ae6ce3a2a280cae30082ef68ede7a1a3efa40),
      .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
     
      // The next set of INITP_xx are for the parity bits
      .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
      
      // The next set of INITP_xx are valid when configured as 36Kb
      .INITP_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_0F(256'h0000000000000000000000000000000000000000000000000000000000000000)
   ) BRAM_TDP_MACRO_inst (
      .DOA(sram_datai),       // Output port-A data, width defined by READ_WIDTH_A parameter
      .DOB(lut_data),       // Output port-B data, width defined by READ_WIDTH_B parameter
      .ADDRA(sram_addr),   // Input port-A address, width defined by Port A depth
      .ADDRB(lut_addr),   // Input port-B address, width defined by Port B depth
      .CLKA(clk),     // 1-bit input port-A clock
      .CLKB(clk),     // 1-bit input port-B clock
      .DIA(sram_datao),       // Input port-A data, width defined by WRITE_WIDTH_A parameter
      .DIB(8'h00),       // Input port-B data, width defined by WRITE_WIDTH_B parameter
      .ENA(1'b1),       // 1-bit input port-A enable
      .ENB(1'b1),       // 1-bit input port-B enable
      .REGCEA(1'b1), // 1-bit input port-A output register enable
      .REGCEB(1'b1), // 1-bit input port-B output register enable
      .RSTA(rst),     // 1-bit input port-A reset
      .RSTB(rst),     // 1-bit input port-B reset
      .WEA({sram_we, sram_we, sram_we, sram_we}),       // Input port-A write enable, width defined by Port A depth
      .WEB(1'b0)        // Input port-B write enable, width defined by Port B depth
   );

   // End of BRAM_TDP_MACRO_inst instantiation

endmodule
